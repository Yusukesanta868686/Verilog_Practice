`define cos1 00000000000000001110110010000011
`define sin1 00000000000000000110000111110111
`define cos2 00000000000000001011010100000100
`define sin2 00000000000000001011010100000100
`define cos3 00000000000000000110000111110111
`define sin3 00000000000000001110110010000011 